drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
drive_router(10'h4, 10'h9, 0);

drive_router(10'h0, 10'h9, 0);
drive_router(10'h1, 10'h5, 0);
drive_router(10'h2, 10'hf, 0);
drive_router(10'h3, 10'h5, 0);
//drive_router(10'h4, 10'h9, 0);

